/**
 * internal_defines.vh
 *
 * This contains the definitions of constants and types that are used by the
 * conFFTi music synthesizer
 **/

`ifndef INTERNAL_DEFINES_VH_
`define INTERNAL_DEFINES_VH_

parameter BAUD_RATE = 31250;
parameter CLOCK_RATE = 50000000;
parameter SAMPLE_RATE = 1600;


`endif  /* INTERNAL_DEFINES_VH_ */