`ifndef OSCILLATOR_VH_
`define OSCILLATOR_VH_

package OSCILLATOR;

typedef enum logic {
  FRONT = 1'b0,
  BACK  = 1'b1
} oscillator_state_t;

endpackage : OSCILLATOR

`endif  /* OSCILLATOR_VH_ */

