module conFFTi (
    input logic clock_50000000,
    input logic clock_184,
    input logic midi_in,
    output logic mixer_out
);

endmodule